library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use IEEE.STD_LOGIC_SIGNED.all;
use IEEE.STD_LOGIC_ARITH.all;
use ieee.numeric_std.all;

-- use IEEE.NUMERIC_STD_UNSIGNED.all;
entity testbench2 is
end;

